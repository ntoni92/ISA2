LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY CARRY_UNIT IS
	GENERIC(N: INTEGER := 9);
	PORT(
		G: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		P: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		c0: IN STD_LOGIC;
		carry: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)	
	);
END ENTITY;

ARCHITECTURE struct OF CARRY_UNIT IS
BEGIN
	carry_gen: FOR i IN 0 TO N-1 GENERATE
		carry(i) <= G(i) OR (c0 AND P(i));
	END GENERATE;
END ARCHITECTURE;