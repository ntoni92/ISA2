jdsvnia
